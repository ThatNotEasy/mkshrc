version https://git-lfs.github.com/spec/v1
oid sha256:7e12d29ab3b59aa86ac0938c2dd97d67f6f14c513c716d3f454e2a2f56c4e423
size 27795
